`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/03/30 20:55:29
// Design Name: 
// Module Name: SCCB
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module top_sccb (
    input  logic clk,
    input  logic reset,
    input  logic btn,
    output logic scl,
    output logic sda
);

    logic [7:0] rom_addr;
    logic [15:0] rom_data;
    logic btn_tick;

    btn_detector U_Btn_Detector (
        .clk(clk),
        .rst(reset),
        .btn(btn),
        .rising_edge_detect(btn_tick),
        .falling_edge_detect(),
        .both_edge_detect()
    );

    SCCB U_SCCB (
        .clk_100MHz(clk),  // 250 count => 400kHz
        .reset(reset),
        .btn_tick(btn_tick),
        .reg_addr(rom_data[15:8]),
        .data(rom_data[7:0]),
        .rom_addr(rom_addr),
        .scl(scl),
        .sda(sda)
    );


    OV7670_config_rom U_ROM (
        .clk (clk),
        .addr(rom_addr),
        .dout(rom_data)
    );
endmodule

module SCCB (
    input logic clk_100MHz,  // 250 count => 400kHz
    input logic reset,
    input logic btn_tick,
    input logic [7:0] reg_addr,
    input logic [7:0] data,
    output logic [7:0] rom_addr,
    output logic scl,
    output logic sda
);

    logic [7:0] counter;
    logic tick_400kHz;

    always_ff @(posedge clk_100MHz, posedge reset) begin
        if (reset) begin
            tick_400kHz <= 0;
            counter <= 0;
        end else begin
            if (counter == 249) begin
                counter <= 0;
                tick_400kHz <= 1'b1;
            end else begin
                counter <= counter + 1;
                tick_400kHz <= 1'b0;
            end
        end
    end

    typedef enum {
        IDLE,
        START,
        DATA,
        STOP,
        CYCLE,
        STAY
    } state_e;

    state_e state;
    logic [1:0] tick_cnt;  // 0, 1, 2, 3
    logic [3:0] bit_cnt;  // 0~15
    logic [1:0] cycle_cnt;  // 0, 1, 2
    logic [7:0] rom_addr_cnt;  // 0~74
    logic [1:0] wait_5us;  // 0, 1
    logic [7:0] id;  // 0x42
    logic start;
    logic [6:0] wait_250us;

    always_ff @(posedge clk_100MHz, posedge reset) begin
        if (reset) begin
            start <= 1'b0;
        end else begin
            if (btn_tick == 1'b1) begin
                start <= 1'b1;
            end else if (tick_400kHz == 1'b1) begin
                start <= 1'b0;
            end
        end
    end

    assign rom_addr = rom_addr_cnt;

    always_comb begin
        scl = 1'b1;
        case(tick_cnt)
        2'b00 : scl = 1'b0; 
        2'b01 : scl = 1'b1;
        2'b10 : scl = 1'b1;
        2'b11 : scl = 1'b0;
        endcase
    end


    always_ff @( posedge clk_100MHz, posedge reset ) begin 
        if(reset)begin
            state <= IDLE;
            wait_5us <= 0;
            tick_cnt <= 1;
            id <= 8'h42;
            cycle_cnt <= 0;
            sda <= 1'b1;
            bit_cnt <= 0;
            rom_addr_cnt <= 0;
            wait_250us <= 0;
        end
        else begin
            case(state)
            IDLE : begin
                rom_addr_cnt <= 0;
                tick_cnt <= 1;
                sda <= 1'b1;
                if(btn_tick)begin
                    state <= START;
                end
                else begin
                    state <= IDLE;
                end
            end

            START : begin
                sda <= 1'b0;
                if(tick_400kHz)begin
                    if(wait_5us == 1)begin
                        wait_5us <= wait_5us + 1;
                        tick_cnt <= 3;
                    end
                    else if(wait_5us == 2)begin
                        state <= DATA;
                        tick_cnt <= 0;
                        wait_5us <= 0;
                        bit_cnt <= 1;
                    end
                    else begin
                        wait_5us <= wait_5us + 1;
                    end
                end
            end

            DATA : begin
                if(tick_400kHz)begin
                    tick_cnt <= tick_cnt + 1;
                    if(tick_cnt == 3)begin
                        if(bit_cnt == 8)begin
                            cycle_cnt <= cycle_cnt + 1;
                            bit_cnt <= 0;
                            sda = 1'b0;
                        end
                        else if(cycle_cnt == 3)begin
                            state <= STOP;
                        end
                        else begin
                            bit_cnt <= bit_cnt + 1;
                            case(cycle_cnt)
                            2'b00 : sda <= id[7-bit_cnt]; 
                            2'b01 : sda <= reg_addr[7-bit_cnt];
                            2'b10 : sda <= data[7-bit_cnt];
                            2'b11 : sda <= 1'b0;
                            endcase
                        end
                    end
                end
            end

            STOP : begin
                cycle_cnt <= 0;
                bit_cnt <= 0;
                if(tick_400kHz)begin
                    if(wait_5us == 1)begin
                        state <= STAY;
                        wait_5us <= 0;
                        sda <= 1'b0;
                    end
                    else begin
                        state <= STOP;
                        wait_5us <= wait_5us + 1;
                        tick_cnt <= 1;
                        sda <= 1'b0;
                    end
                end
            end

            STAY : begin
                sda <= 1'b1;
                if(rom_addr_cnt == 74)begin
                    state <= IDLE;
                end
                else begin
                    if(tick_400kHz)begin
                        if(wait_250us == 99)begin
                            state <= START;
                            rom_addr_cnt <= rom_addr_cnt + 1;
                            wait_250us <= 0;
                        end
                        else begin
                            state <= STAY;
                            wait_250us <= wait_250us + 1;
                        end
                    end
                end
            end
            endcase
        end
    end

endmodule

module OV7670_config_rom (
    input logic clk,
    input logic [7:0] addr,
    output logic [15:0] dout
);

    //FFFF is end of rom, FFF0 is delay
    always @(posedge clk) begin
        case (addr)
            0: dout <= 16'h12_80;  //reset
            1: dout <= 16'hFF_F0;  //delay
            2:
            dout <= 16'h12_14;  // COM7,     set RGB color output and set QVGA
            3: dout <= 16'h11_80;  // CLKRC     internal PLL matches input clock
            4: dout <= 16'h0C_04;  // COM3,     default settings
            5: dout <= 16'h3E_19;  // COM14,    no scaling, normal pclock
            6: dout <= 16'h04_00;  // COM1,     disable CCIR656
            7: dout <= 16'h40_d0;  //COM15,     RGB565, full output range
            8: dout <= 16'h3a_04;  //TSLB       
            9: dout <= 16'h14_18;  //COM9       MAX AGC value x4
            10: dout <= 16'h4F_B3;  //MTX1       
            11: dout <= 16'h50_B3;  //MTX2
            12: dout <= 16'h51_00;  //MTX3
            13: dout <= 16'h52_3d;  //MTX4
            14: dout <= 16'h53_A7;  //MTX5
            15: dout <= 16'h54_E4;  //MTX6
            16: dout <= 16'h58_9E;  //MTXS
            17:
            dout <= 16'h3D_C0; //COM13      sets gamma enable, does not preserve reserved bits, may be wrong?
            18: dout <= 16'h17_15;  //HSTART     start high 8 bits 
            19:
            dout <= 16'h18_03; //HSTOP      stop high 8 bits //these kill the odd colored line
            20: dout <= 16'h32_00;  //91  //HREF       edge offset
            21: dout <= 16'h19_03;  //VSTART     start high 8 bits
            22: dout <= 16'h1A_7B;  //VSTOP      stop high 8 bits
            23: dout <= 16'h03_00;  // 00 //VREF       vsync edge offset
            24: dout <= 16'h0F_41;  //COM6       reset timings
            25:
            dout <= 16'h1E_00; //MVFP       disable mirror / flip //might have magic value of 03
            26: dout <= 16'h33_0B;  //CHLF       //magic value from the internet
            27: dout <= 16'h3C_78;  //COM12      no HREF when VSYNC low
            28: dout <= 16'h69_00;  //GFIX       fix gain control
            29: dout <= 16'h74_00;  //REG74      Digital gain control
            30:
            dout <= 16'hB0_84; //RSVD       magic value from the internet *required* for good color
            31: dout <= 16'hB1_0c;  //ABLC1
            32: dout <= 16'hB2_0e;  //RSVD       more magic internet values
            33: dout <= 16'hB3_80;  //THL_ST
            //begin mystery scaling numbers
            34: dout <= 16'h70_3a;
            35: dout <= 16'h71_35;
            36: dout <= 16'h72_11;
            37: dout <= 16'h73_f1;
            38: dout <= 16'ha2_02;
            //gamma curve values
            39: dout <= 16'h7a_20;
            40: dout <= 16'h7b_10;
            41: dout <= 16'h7c_1e;
            42: dout <= 16'h7d_35;
            43: dout <= 16'h7e_5a;
            44: dout <= 16'h7f_69;
            45: dout <= 16'h80_76;
            46: dout <= 16'h81_80;
            47: dout <= 16'h82_88;
            48: dout <= 16'h83_8f;
            49: dout <= 16'h84_96;
            50: dout <= 16'h85_a3;
            51: dout <= 16'h86_af;
            52: dout <= 16'h87_c4;
            53: dout <= 16'h88_d7;
            54: dout <= 16'h89_e8;
            //AGC and AEC
            55: dout <= 16'h13_e0;  //COM8, disable AGC / AEC
            56: dout <= 16'h00_00;  //set gain reg to 0 for AGC
            57: dout <= 16'h10_00;  //set ARCJ reg to 0
            58: dout <= 16'h0d_40;  //magic reserved bit for COM4
            59: dout <= 16'h14_18;  //COM9, 4x gain + magic bit
            60: dout <= 16'ha5_05;  // BD50MAX
            61: dout <= 16'hab_07;  //DB60MAX
            62: dout <= 16'h24_95;  //AGC upper limit
            63: dout <= 16'h25_33;  //AGC lower limit
            64: dout <= 16'h26_e3;  //AGC/AEC fast mode op region
            65: dout <= 16'h9f_78;  //HAECC1
            66: dout <= 16'ha0_68;  //HAECC2
            67: dout <= 16'ha1_03;  //magic
            68: dout <= 16'ha6_d8;  //HAECC3
            69: dout <= 16'ha7_d8;  //HAECC4
            70: dout <= 16'ha8_f0;  //HAECC5
            71: dout <= 16'ha9_90;  //HAECC6
            72: dout <= 16'haa_94;  //HAECC7
            73: dout <= 16'h13_e7;  //COM8, enable AGC / AEC
            74: dout <= 16'h69_07;
            default: dout <= 16'hFF_FF;  //mark end of ROM
        endcase
    end
endmodule

// module btn_detector (
//     input  logic clk,
//     input  logic reset,
//     input  logic btn,
//     output logic rising_edge,
//     output logic falling_edge,
//     output logic both_edge
// );

//     reg [3:0] shift_reg;
//     reg q_reg;
//     reg [$clog2(100_000)-1:0] tick_cnt;
//     reg tick;
//     wire debounce;

//     always @(posedge clk, posedge reset) begin
//         if (reset) begin
//             tick_cnt <= 0;
//             tick <= 0;
//         end else begin
//             if (tick_cnt <= 100_000 - 1) begin
//                 tick_cnt <= 0;
//                 tick <= 1'b1;
//             end else begin
//                 tick_cnt <= tick_cnt + 1;
//                 tick <= 1'b0;
//             end
//         end
//     end

//     always @(posedge clk, posedge reset) begin
//         if (reset) begin
//             shift_reg <= 0;
//         end else begin
//             if (tick) begin
//                 shift_reg <= {
//                     btn, shift_reg[3:1]
//                 };  // shift_reg = shift_reg >> 1;
//                 // shift_reg <= {shift_reg[2:0], in};  // shift_reg = shift_reg << 1;
//             end
//         end
//     end

//     assign debounce = &shift_reg; // shift_reg[3] & shift_reg[2] & shift_reg[1] & shift_reg[0]

//     always @(posedge clk, posedge reset) begin
//         if (reset) begin
//             q_reg <= 1'b0;
//         end else begin
//             q_reg <= debounce;
//         end
//     end

//     assign rising_edge = debounce & ~q_reg;
//     assign falling_edge = ~debounce & q_reg;
//     assign both_edge = rising_edge | falling_edge;

// endmodule





