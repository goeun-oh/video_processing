`timescale 1ns/1ps


module SCCB_Controller(
    input logic clk,
    input logic reset,
    output logic scl,
    output logic sda
);
    typedef enum  { IDLE,  } name;

endmodule