
module font_rom (
    input  logic [6:0] char_code,   // ASCII 코드 (0~127)
    input  logic [2:0] row_index,   // 글자 한 줄 (0~7)
    output logic [7:0] row_data     // 출력: 해당 줄의 비트맵
);
    // 글자 비트맵 ROM [ASCII][Row]
    logic [7:0] font [0:127][0:7];

    initial begin
        // 'G'
        font["G"][0] = 8'b00111110;
        font["G"][1] = 8'b01100000;
        font["G"][2] = 8'b11000000;
        font["G"][3] = 8'b11001110;
        font["G"][4] = 8'b11000010;
        font["G"][5] = 8'b01100010;
        font["G"][6] = 8'b00111100;
        font["G"][7] = 8'b00000000;

        // 'A'
        font["A"][0] = 8'b00011000;
        font["A"][1] = 8'b00100100;
        font["A"][2] = 8'b01000010;
        font["A"][3] = 8'b01000010;
        font["A"][4] = 8'b01111110;
        font["A"][5] = 8'b01000010;
        font["A"][6] = 8'b01000010;
        font["A"][7] = 8'b00000000;

        // 'M'
        font["M"][0] = 8'b10000001;
        font["M"][1] = 8'b11000011;
        font["M"][2] = 8'b10100101;
        font["M"][3] = 8'b10011001;
        font["M"][4] = 8'b10000001;
        font["M"][5] = 8'b10000001;
        font["M"][6] = 8'b10000001;
        font["M"][7] = 8'b00000000;

        // 'E'
        font["E"][0] = 8'b01111110;
        font["E"][1] = 8'b01000000;
        font["E"][2] = 8'b01111000;
        font["E"][3] = 8'b01000000;
        font["E"][4] = 8'b01000000;
        font["E"][5] = 8'b01111110;
        font["E"][6] = 8'b00000000;
        font["E"][7] = 8'b00000000;

        // 'O'
        font["O"][0] = 8'b00111100;
        font["O"][1] = 8'b01000010;
        font["O"][2] = 8'b10000001;
        font["O"][3] = 8'b10000001;
        font["O"][4] = 8'b10000001;
        font["O"][5] = 8'b01000010;
        font["O"][6] = 8'b00111100;
        font["O"][7] = 8'b00000000;

        // 'V'
        font["V"][0] = 8'b10000001;
        font["V"][1] = 8'b10000001;
        font["V"][2] = 8'b01000010;
        font["V"][3] = 8'b01000010;
        font["V"][4] = 8'b00100100;
        font["V"][5] = 8'b00011000;
        font["V"][6] = 8'b00011000;
        font["V"][7] = 8'b00000000;

        // 'R'
        font["R"][0] = 8'b01111110;
        font["R"][1] = 8'b01000010;
        font["R"][2] = 8'b01111110;
        font["R"][3] = 8'b01001000;
        font["R"][4] = 8'b01000100;
        font["R"][5] = 8'b01000010;
        font["R"][6] = 8'b00000000;
        font["R"][7] = 8'b00000000;

        // ' ' (space)
        font[" "][0] = 8'b00000000;
        font[" "][1] = 8'b00000000;
        font[" "][2] = 8'b00000000;
        font[" "][3] = 8'b00000000;
        font[" "][4] = 8'b00000000;
        font[" "][5] = 8'b00000000;
        font[" "][6] = 8'b00000000;
        font[" "][7] = 8'b00000000;
    end

    assign row_data = font[char_code][row_index];
endmodule
